// Примеры использования см. в конце кода

// Главное правило:
// "Нельзя использовать BRAM только для записи без последующего чтения и использования результата.
// В ПЛИС всё, что не влияет на выходы, удаляется."
// Поэтому даже в «режиме записи» вы обязаны прочитать и отобразить/вывести данные — тогда синтезатор поймёт, что BRAM нужен.

module bram_rw_controller
(
    input        clk,

    // Интерфейс записи
    input        wr_en,
    input  [3:0] wr_addr,
    input  [7:0] wr_data,

    // Интерфейс чтения
    input        rd_en,
    input  [3:0] rd_addr,
    output reg [7:0] rd_data
);

// ================================================================================
wire [7:0] bram_dout;         // выход BRAM
wire       bram_ce;           // разрешение работы порта
wire       bram_oce;          // разрешение вывода данных
wire       bram_wre;          // разрешение записи
wire [3:0] bram_ad;           // адрес (общий для чтения и записи)

// ================================================================================

// Порт активен, если есть запрос на чтение ИЛИ запись
assign bram_ce  = rd_en | wr_en;

// Запись разрешена ТОЛЬКО при wr_en (и не при одновременном rd_en!)
// В SP-режиме одновременная запись и чтение — неопределённое поведение!
// Поэтому приоритет: запись, если wr_en = 1; иначе — чтение.
assign bram_wre = wr_en;
assign bram_ad  = wr_en ? wr_addr : rd_addr;

// Выход разрешён ТОЛЬКО при чтении (и отсутствии записи в тот же такт)
// (на практике: если wr_en = 1, чтение в этот такт игнорируется)
assign bram_oce = rd_en & (~wr_en);

// ================================================================================

bram_sp_init bram_inst (
    .dout(bram_dout),
    .clk(clk),
    .oce(bram_oce),
    .ce(bram_ce),
    .reset(1'b0),       // сброс не используется — память инициализирована
    .wre(bram_wre),
    .ad(bram_ad),
    .din(wr_data)       // при записи — wr_data, при чтении — безразлично
);

// ================================================================================

// ----------------------------------------------------------------------
// Регистрация выходных данных (registered read)
// rd_data обновляется на следующем такте после rd_en
// ----------------------------------------------------------------------
always @(posedge clk) begin
    if (rd_en && !wr_en)  // читаем только если не пишем в тот же такт
        rd_data <= bram_dout;
end

endmodule



// ПРИМЕРЫ ИСПОЛЬЗОВАНИЯ

// 1. только для чтения
    //bram_rw_controller bram_inst (
    //    .clk(clk),
    //    .wr_en(1'b0),           // запись отключена
    //    .wr_addr(3'd0),
    //    .wr_data(8'd0),
    //    .rd_en(rd_en),
    //    .rd_addr(addr),
    //    .rd_data(rd_data)
    //);

// 2. только для записи
    //bram_rw_controller bram_inst (
    //    .clk(clk),
    //    .wr_en(wr_en),
    //    .wr_addr(addr),          // пишем в адрес 0
    //    .wr_data(data_to_write),
    //    .rd_en(rd_en),
    //    .rd_addr(addr),          // читаем тот же адрес
    //    .rd_data(rd_data)
    //);

// 3. чтение + запись
    //bram_rw u_bram (
    //    .clk(clk),
    //    .wr_en(wr_en),
    //    .wr_addr(wr_addr),
    //    .wr_data(wr_data),
    //    .rd_en(rd_en),
    //    .rd_addr(rd_addr),
    //    .rd_data(rd_data)
    //);
